*##########################################################################################
* Copyright (c) 2023 Dolphin Technology, Inc.
* This netlist is proprietary and confidential information of
* Dolphin Technology, Inc. and can only be used or viewed
* under license or with written permission from Dolphin Technology, Inc.
*##########################################################################################
* /data/projects/stdcells/scripts_svn_update_flow/Update_property_flow/lvsNetlist.pl -c dti_55g_10t_nor2x1 -p /data/projects/stdcells/scripts_svn_update_flow/Update_property_flow/params/params55.sp -s netlist -d lvs -nglob
* dt35-linux:/data/projects/stdcells/REPOSITORY_RV003/ckt/tsmc55 
* dti_55g_10t_nor2x1.ckt generated on 6/5/2023 at 10:3:45
*##########################################################################################
* Dependencies
*##########################################################################################

.param wnd=1u wpd=1u

.option scale=1

.global vdd vss vddps vddcs
* DAMN, don't know where the cell is 
.subckt dti_55g_10t_nor2x1 VDD VSS A B Z
mp1 Z A N1N71 VDD pch l=0.06u w=0.735u
mn1 Z A VSS VSS nch l=0.06u w=0.525u
mn2 Z B VSS VSS nch l=0.06u w=0.525u
mp2 N1N71 B VDD VDD pch l=0.06u w=0.735u
.ends

