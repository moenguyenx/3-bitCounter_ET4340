*##########################################################################################
* Copyright (c) 2023 Dolphin Technology, Inc.
* This netlist is proprietary and confidential information of
* Dolphin Technology, Inc. and can only be used or viewed
* under license or with written permission from Dolphin Technology, Inc.
*##########################################################################################
* /data/projects/stdcells/scripts_svn_update_flow/Update_property_flow/lvsNetlist.pl -c dti_55g_10t_or2x1 -p /data/projects/stdcells/scripts_svn_update_flow/Update_property_flow/params/params55.sp -s netlist -d lvs -nglob
* dt35-linux:/data/projects/stdcells/REPOSITORY_RV003/ckt/tsmc55 
* dti_55g_10t_or2x1.ckt generated on 6/5/2023 at 11:0:11
*##########################################################################################
* Dependencies
*##########################################################################################

.param wnd=1u wpd=1u

.option scale=1

.global vdd vss vddps vddcs
* DAMN, don't know where the cell is 
.subckt dti_55g_10t_or2x1 VDD VSS Z A B
mp2 N1N47 A N1N71 VDD pch l=0.06u w=0.735u
mp1 Z N1N47 VDD VDD pch l=0.06u w=0.735u
mn1 Z N1N47 VSS VSS nch l=0.06u w=0.525u
mn2 N1N47 A VSS VSS nch l=0.06u w=0.525u
mp3 N1N71 B VDD VDD pch l=0.06u w=0.735u
mn3 N1N47 B VSS VSS nch l=0.06u w=0.525u
.ends

