*##########################################################################################
* Copyright (c) 2023 Dolphin Technology, Inc.
* This netlist is proprietary and confidential information of
* Dolphin Technology, Inc. and can only be used or viewed
* under license or with written permission from Dolphin Technology, Inc.
*##########################################################################################
* /data/projects/stdcells/scripts_svn_update_flow/Update_property_flow/lvsNetlist.pl -c dti_55g_10t_xor2x1 -p /data/projects/stdcells/scripts_svn_update_flow/Update_property_flow/params/params55.sp -s netlist -d lvs -nglob
* dt35-linux:/data/projects/stdcells/REPOSITORY_RV003/ckt/tsmc55 
* dti_55g_10t_xor2x1.ckt generated on 6/5/2023 at 16:38:32
*##########################################################################################
* Dependencies
*##########################################################################################

.param wnd=1u wpd=1u

.option scale=1

.global vdd vss vddps vddcs
* DAMN, don't know where the cell is 
.subckt dti_55g_10t_xor2x1 VDD VSS B Z A
x1i55 VDD VSS A N1N56 dti_gen_inv wn=0.525u wp=0.525u
x1i62 VDD VSS N1N56 N1N58 dti_gen_inv wn=0.525u wp=0.525u
x1i57 VDD VSS N1N27 Z dti_gen_inv wn=0.525u wp=0.525u
x1i63 VDD VSS B N1N23 dti_gen_inv wn=0.525u wp=0.525u
x1i61 VDD VSS N1N23 B N1N58 N1N27 dti_gen_tx wn=0.525u wp=0.525u
x1i15 VDD VSS B N1N23 N1N56 N1N27 dti_gen_tx wn=0.525u wp=0.525u
.ends

* DAMN, don't know where the cell is 
.subckt dti_gen_inv VDD VSS A Z ln=0.06u lp=0.06u wn=0.15u wp=0.15u
m1i3 Z A VDD VDD pch l=lp w=wp
m1i4 Z A VSS VSS nch l=ln w=wn
.ends

* DAMN, don't know where the cell is 
.subckt dti_gen_tx VDD VSS PG NG IN OUT wn=0.15u wp=0.15u
m1i3 IN PG OUT VDD pch l=0.06u w=wp
m1i2 IN NG OUT VSS nch l=0.06u w=wn
.ends

