*##########################################################################################
* Copyright (c) 2023 Dolphin Technology, Inc.
* This netlist is proprietary and confidential information of
* Dolphin Technology, Inc. and can only be used or viewed
* under license or with written permission from Dolphin Technology, Inc.
*##########################################################################################
* /data/projects/stdcells/scripts_svn_update_flow/Update_property_flow/lvsNetlist.pl -c dti_55g_10t_and3x1 -p /data/projects/stdcells/scripts_svn_update_flow/Update_property_flow/params/params55.sp -s netlist -d lvs -nglob
* dt35-linux:/data/projects/stdcells/REPOSITORY_RV003/ckt/tsmc55 
* dti_55g_10t_and3x1.ckt generated on 6/2/2023 at 17:22:35
*##########################################################################################
* Dependencies
*##########################################################################################

.param wnd=1u wpd=1u

.option scale=1

.global vdd vss vddps vddcs
* DAMN, don't know where the cell is 
.subckt dti_55g_10t_and3x1 VDD VSS C Z A B
mp4 N1N47 C VDD VDD pch l=0.06u w=0.735u
mp2 N1N47 A VDD VDD pch l=0.06u w=0.735u
mp1 Z N1N47 VDD VDD pch l=0.06u w=0.735u
mn1 Z N1N47 VSS VSS nch l=0.06u w=0.525u
mp3 N1N47 B VDD VDD pch l=0.06u w=0.735u
mn2 N1N47 A N1N43 VSS nch l=0.06u w=0.525u
mn3 N1N43 B N1N71 VSS nch l=0.06u w=0.525u
mn4 N1N71 C VSS VSS nch l=0.06u w=0.525u
.ends

